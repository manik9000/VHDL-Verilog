
library ieee
